// Intersection controller module

module intersectionController
(
	input [5:0] perTime, 
	input [5:0] handTime, 
	input [5:0] redTime, 
	input [5:0] yellowTime, 
	input [5:0] greenTime,

	output fsmPedControl, 
	output fsmCarControl
);

// Module definitions


endmodule