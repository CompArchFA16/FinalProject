// 2Hz blink timer module

module blinkTimer
(
	input clk,
	input reset,
	output blink
);

wire [14:0] upCounter;

always @(posedge clk)

	// Up counter
	if (reset) begin
		upCounter <= 8'b0 ;
	end else if (enable) begin
		upCounter <= upCounter + 1;
	end

	assign blink = &upCounter;

endmodule