// Intersection controller module

module intersectionController
(
	// Def
);

endmodule